`timescale 1ns / 1ps

module Decoder_TB(

    );
endmodule
